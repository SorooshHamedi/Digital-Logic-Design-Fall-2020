`timescale 1ns/1ns
module nBitInverter(A, w);
	parameter SIZE = 8;
	input [SIZE-1:0]A;
	output [SIZE-1:0]w;

	genvar i;
	generate
		for(i=0; i<SIZE; i=i+1) begin: inverter
			assign #(5,7) w[i] = ~A[i];
		end
	endgenerate
endmodule
