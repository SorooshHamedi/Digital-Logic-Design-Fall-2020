`timescale 1ns/1ns
module nBitAdder(A, B, sum, carryOut);
	parameter SIZE = 8;
	input [SIZE-1:0]A, B;
	output [SIZE-1:0]sum;
	output carryOut;
	wire [SIZE/2:0]carry;
	
	assign carry[0] = 1'b0;
	assign carryOut = carry[SIZE/2];

	genvar i;
	generate
		for(i=0; i<SIZE/2; i=i+1) begin
			TwoBitMuxBasedAdder tma(.A({A[i*2+1], A[i*2]}), .B({B[i*2+1], B[i*2]}), .carryIn(carry[i]), .sum({sum[i*2+1], sum[i*2]}), .carryOut(carry[i+1]));
		end
	endgenerate
endmodule
	