`timescale 1ns/1ns
module BufIf0(input A, input en, output w);
	bufif0 #(17,19,19) buff(w,A,en);
endmodule
